library verilog;
use verilog.vl_types.all;
entity processor is
end processor;
